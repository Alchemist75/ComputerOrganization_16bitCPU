----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:40:11 12/05/2017 
-- Design Name: 
-- Module Name:    RstController - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RstController is
    Port ( rst : in  STD_LOGIC;
           FLASH_FINISH : in  STD_LOGIC;
           rst_out : out  STD_LOGIC);
end RstController;

architecture Behavioral of RstController is

begin

	rst_out <= rst and FLASH_FINISH;

end Behavioral;

